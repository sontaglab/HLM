module rca2 ();
//-------------Input Ports Declarations-----------------------------
input;
//-------------Output Ports Declarations-----------------------------
output s;
assign s = ;
endmodule