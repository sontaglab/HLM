module rca2 (x_1,x_2,x_3,x_4,s);
//-------------Input Ports Declarations-----------------------------
input x_1,x_2,x_3,x_4;
//-------------Output Ports Declarations-----------------------------
output s;
//-------------Logic-----------------------------------------------
assign s =  ( ~x_1 & ~x_2 & ~x_3 & ~x_4 ) | ( ~x_1 & ~x_2 & ~x_3 & x_4 ) | ( ~x_1 & ~x_2 & x_3 & ~x_4 ) | ( ~x_1 & x_2 & x_3 & ~x_4 ) | ( x_1 & ~x_2 & ~x_3 & ~x_4 ) | ( x_1 & ~x_2 & x_3 & ~x_4 ) | ( x_1 & x_2 & ~x_3 & ~x_4 ) | ( x_1 & x_2 & ~x_3 & x_4 ) | ( x_1 & x_2 & x_3 & ~x_4 ) | ( x_1 & x_2 & x_3 & x_4 );
endmodule